
module mycore
(
	input         clk,
	input         reset
	

);


endmodule
