//-------------------------------------------------------------------------------------------------
module rom
//-------------------------------------------------------------------------------------------------
#
(
	parameter DW = 8,
	parameter AW = 14,
	parameter FN = ""
)
(
	input  wire          clock,
	input  wire          ce,

	output reg  [DW-1:0] data_out,
	output reg  [AW-1:0] out_address
);
//-------------------------------------------------------------------------------------------------

reg[DW-1:0] d[(2**AW)-1:0];
initial $readmemh(FN, d, 0);

always @(posedge clock) begin
	if(ce) 
	begin
		out_address <= out_address + 1'd1;		
		data_out <= d[out_address];		
	end
end

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
