//-------------------------------------------------------------------------------------------------
module rommif
//-------------------------------------------------------------------------------------------------
#
(
	parameter DW = 8,
	parameter AW = 14,
	parameter FN = ""
)
(
	input  wire            clock,
	input  wire            ce,
	input  wire  [AW-1:0]  in_address,

	output reg   [DW-1:0]  data_out
);

//-------------------------------------------------------------------------------------------------

reg[DW-1:0] d[(2**AW)-1:0];
initial $readmemb(FN, d, 0);

always @(posedge clock) begin
	data_out <= d[in_address];	
end

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
